
`define RADD            4'b0010    // Signed addition (A + B)
`define MUL_ALU         4'b1100
`define LSW             4'b0110  
`define RB              4'b0001    // Pass-through B (Output = B)
`define LDR             4'b1001  
`define RSUB            4'b0011    // Signed subtraction (A - B)
`define LDSW_FULL_ALU   4'b1000   
`define MOVSW_ALU       4'b1010



