module rom #(
    parameter WIDTH = 8,
    parameter DEPTH = 256,
    parameter ADDR_WIDTH = 8
) (
    input logic clk,
    input logic [ADDR_WIDTH-1:0] addr,
    output logic [WIDTH-1:0] dout
);
    logic [WIDTH-1:0] memory [0:DEPTH-1];

    assign dout = memory[addr];  // Combinational read

    initial begin
        // Noisy samples at 0-255
        memory[0]   = 8'hF6;
        memory[1]   = 8'h02;
        memory[2]   = 8'h0F;
        memory[3]   = 8'h1A;
        memory[4]   = 8'h10;
        memory[5]   = 8'h13;
        memory[6]   = 8'h2A;
        memory[7]   = 8'h1F;
        memory[8]   = 8'h2C;
        memory[9]   = 8'h2C;
        memory[10]  = 8'h3B;
        memory[11]  = 8'h2D;
        memory[12]  = 8'h2F;
        memory[13]  = 8'h43;
        memory[14]  = 8'h3C;
        memory[15]  = 8'h50;
        memory[16]  = 8'h4F;
        memory[17]  = 8'h40;
        memory[18]  = 8'h55;
        memory[19]  = 8'h4A;
        memory[20]  = 8'h61;
        memory[21]  = 8'h53;
        memory[22]  = 8'h61;
        memory[23]  = 8'h57;
        memory[24]  = 8'h5D;
        memory[25]  = 8'h61;
        memory[26]  = 8'h6D;
        memory[27]  = 8'h70;
        memory[28]  = 8'h62;
        memory[29]  = 8'h69;
        memory[30]  = 8'h65;
        memory[31]  = 8'h5E;
        memory[32]  = 8'h73;
        memory[33]  = 8'h68;
        memory[34]  = 8'h5D;
        memory[35]  = 8'h65;
        memory[36]  = 8'h62;
        memory[37]  = 8'h65;
        memory[38]  = 8'h55;
        memory[39]  = 8'h5F;
        memory[40]  = 8'h53;
        memory[41]  = 8'h58;
        memory[42]  = 8'h51;
        memory[43]  = 8'h4F;
        memory[44]  = 8'h58;
        memory[45]  = 8'h5D;
        memory[46]  = 8'h48;
        memory[47]  = 8'h45;
        memory[48]  = 8'h41;
        memory[49]  = 8'h50;
        memory[50]  = 8'h49;
        memory[51]  = 8'h3A;
        memory[52]  = 8'h2C;
        memory[53]  = 8'h3C;
        memory[54]  = 8'h28;
        memory[55]  = 8'h30;
        memory[56]  = 8'h31;
        memory[57]  = 8'h1A;
        memory[58]  = 8'h13;
        memory[59]  = 8'h13;
        memory[60]  = 8'h0B;
        memory[61]  = 8'h04;
        memory[62]  = 8'h10;
        memory[63]  = 8'h09;
        memory[64]  = 8'h06;
        memory[65]  = 8'h02;
        memory[66]  = 8'hED;
        memory[67]  = 8'hEA;
        memory[68]  = 8'hE2;
        memory[69]  = 8'hEF;
        memory[70]  = 8'hD6;
        memory[71]  = 8'hD5;
        memory[72]  = 8'hDC;
        memory[73]  = 8'hDB;
        memory[74]  = 8'hCB;
        memory[75]  = 8'hCE;
        memory[76]  = 8'hCC;
        memory[77]  = 8'hC1;
        memory[78]  = 8'hB4;
        memory[79]  = 8'hBE;
        memory[80]  = 8'hBD;
        memory[81]  = 8'hB9;
        memory[82]  = 8'hA8;
        memory[83]  = 8'hB6;
        memory[84]  = 8'hB5;
        memory[85]  = 8'h9E;
        memory[86]  = 8'hB1;
        memory[87]  = 8'hA8;
        memory[88]  = 8'hA6;
        memory[89]  = 8'hA1;
        memory[90]  = 8'hAA;
        memory[91]  = 8'hA6;
        memory[92]  = 8'hA5;
        memory[93]  = 8'hA2;
        memory[94]  = 8'h99;
        memory[95]  = 8'h94;
        memory[96]  = 8'h9F;
        memory[97]  = 8'hA0;
        memory[98]  = 8'hA6;
        memory[99]  = 8'hA0;
        memory[100] = 8'hA2;
        memory[101] = 8'hA6;
        memory[102] = 8'hAA;
        memory[103] = 8'h9C;
        memory[104] = 8'hAD;
        memory[105] = 8'hAC;
        memory[106] = 8'hA6;
        memory[107] = 8'hAA;
        memory[108] = 8'hAF;
        memory[109] = 8'hA7;
        memory[110] = 8'hA4;
        memory[111] = 8'hBB;
        memory[112] = 8'hAC;
        memory[113] = 8'hB7;
        memory[114] = 8'hCA;
        memory[115] = 8'hBB;
        memory[116] = 8'hD3;
        memory[117] = 8'hD5;
        memory[118] = 8'hD2;
        memory[119] = 8'hD5;
        memory[120] = 8'hE6;
        memory[121] = 8'hDA;
        memory[122] = 8'hD9;
        memory[123] = 8'hEC;
        memory[124] = 8'hF8;
        memory[125] = 8'hE7;
        memory[126] = 8'hEC;
        memory[127] = 8'hFE;
        memory[128] = 8'h0A;
        memory[129] = 8'hFF;
        memory[130] = 8'h06;
        memory[131] = 8'h08;
        memory[132] = 8'h09;
        memory[133] = 8'h1C;
        memory[134] = 8'h21;
        memory[135] = 8'h2D;
        memory[136] = 8'h1D;
        memory[137] = 8'h2D;
        memory[138] = 8'h33;
        memory[139] = 8'h3F;
        memory[140] = 8'h41;
        memory[141] = 8'h3C;
        memory[142] = 8'h4C;
        memory[143] = 8'h49;
        memory[144] = 8'h48;
        memory[145] = 8'h45;
        memory[146] = 8'h4E;
        memory[147] = 8'h59;
        memory[148] = 8'h54;
        memory[149] = 8'h63;
        memory[150] = 8'h5D;
        memory[151] = 8'h58;
        memory[152] = 8'h65;
        memory[153] = 8'h6C;
        memory[154] = 8'h6D;
        memory[155] = 8'h6D;
        memory[156] = 8'h66;
        memory[157] = 8'h70;
        memory[158] = 8'h5B;
        memory[159] = 8'h5B;
        memory[160] = 8'h6F;
        memory[161] = 8'h71;
        memory[162] = 8'h68;
        memory[163] = 8'h5F;
        memory[164] = 8'h6F;
        memory[165] = 8'h63;
        memory[166] = 8'h6A;
        memory[167] = 8'h5F;
        memory[168] = 8'h58;
        memory[169] = 8'h5B;
        memory[170] = 8'h5D;
        memory[171] = 8'h5C;
        memory[172] = 8'h4E;
        memory[173] = 8'h50;
        memory[174] = 8'h4E;
        memory[175] = 8'h4F;
        memory[176] = 8'h49;
        memory[177] = 8'h4A;
        memory[178] = 8'h48;
        memory[179] = 8'h40;
        memory[180] = 8'h3E;
        memory[181] = 8'h40;
        memory[182] = 8'h2B;
        memory[183] = 8'h2A;
        memory[184] = 8'h24;
        memory[185] = 8'h22;
        memory[186] = 8'h16;
        memory[187] = 8'h24;
        memory[188] = 8'h18;
        memory[189] = 8'h03;
        memory[190] = 8'h11;
        memory[191] = 8'hFC;
        memory[192] = 8'h03;
        memory[193] = 8'hF9;
        memory[194] = 8'h02;
        memory[195] = 8'hF0;
        memory[196] = 8'hF0;
        memory[197] = 8'hF2;
        memory[198] = 8'hEA;
        memory[199] = 8'hD7;
        memory[200] = 8'hDA;
        memory[201] = 8'hCD;
        memory[202] = 8'hC6;
        memory[203] = 8'hD7;
        memory[204] = 8'hC3;
        memory[205] = 8'hBD;
        memory[206] = 8'hBA;
        memory[207] = 8'hB4;
        memory[208] = 8'hC0;
        memory[209] = 8'hC1;
        memory[210] = 8'hAD;
        memory[211] = 8'hAA;
        memory[212] = 8'hB1;
        memory[213] = 8'hA6;
        memory[214] = 8'hB2;
        memory[215] = 8'hA1;
        memory[216] = 8'hA1;
        memory[217] = 8'h99;
        memory[218] = 8'hAB;
        memory[219] = 8'h97;
        memory[220] = 8'h9C;
        memory[221] = 8'hA4;
        memory[222] = 8'h98;
        memory[223] = 8'hA3;
        memory[224] = 8'h8D;
        memory[225] = 8'h97;
        memory[226] = 8'hA1;
        memory[227] = 8'hA0;
        memory[228] = 8'h9C;
        memory[229] = 8'hA1;
        memory[230] = 8'h9E;
        memory[231] = 8'hA1;
        memory[232] = 8'hA3;
        memory[233] = 8'hAF;
        memory[234] = 8'hB1;
        memory[235] = 8'hB2;
        memory[236] = 8'hB4;
        memory[237] = 8'hA2;
        memory[238] = 8'hA9;
        memory[239] = 8'hB0;
        memory[240] = 8'hB1;
        memory[241] = 8'hBA;
        memory[242] = 8'hBE;
        memory[243] = 8'hC4;
        memory[244] = 8'hD1;
        memory[245] = 8'hD2;
        memory[246] = 8'hD9;
        memory[247] = 8'hDC;
        memory[248] = 8'hE2;
        memory[249] = 8'hD1;
        memory[250] = 8'hE5;
        memory[251] = 8'hE0;
        memory[252] = 8'hED;
        memory[253] = 8'hFC;
        memory[254] = 8'hF4;
        memory[255] = 8'hEF;
        
        
    end

  always_comb begin
  $display("ROM: addr=%h, dout=%h, memory[addr]=%h", addr, dout, memory[addr]);
end
endmodule